module tlm;
  
endmodule
