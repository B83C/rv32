`ifndef DEFS_SVH 
`define DEFS_SVH
typedef enum {
  ADD = 0,
  SLL,
  SLT,
  SLTU,
  XOR,
  SRLA,
  OR,
  AND
} alu_op_t;

`endif
