module alu_ctrl #(
  IR_WIDTH = 6'd32
)(
  input [IR_WIDTH - 1: 0] ir��
  output 
);

endmodule
