module mmio;
endmodule
