module mmio(
  input [31:0] addr,
  output addr_mem, 
  output [31:0] data 
);

assign data = 




endmodule
